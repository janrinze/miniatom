/*

  character generator

*/


module charGen (
	input [9:0] address,
	output [7:0]dout);
always @ (address)
begin
case (address)
3 :dout = 8'b00011100 ;
4 :dout = 8'b00100010 ;
5 :dout = 8'b00000010 ;
6 :dout = 8'b00011010 ;
7 :dout = 8'b00101010 ;
8 :dout = 8'b00101010 ;
9 :dout = 8'b00011100 ;
19 :dout = 8'b00001000 ;
20 :dout = 8'b00010100 ;
21 :dout = 8'b00100010 ;
22 :dout = 8'b00100010 ;
23 :dout = 8'b00111110 ;
24 :dout = 8'b00100010 ;
25 :dout = 8'b00100010 ;
35 :dout = 8'b00111100 ;
36 :dout = 8'b00010010 ;
37 :dout = 8'b00010010 ;
38 :dout = 8'b00011100 ;
39 :dout = 8'b00010010 ;
40 :dout = 8'b00010010 ;
41 :dout = 8'b00111100 ;
51 :dout = 8'b00011100 ;
52 :dout = 8'b00100010 ;
53 :dout = 8'b00100000 ;
54 :dout = 8'b00100000 ;
55 :dout = 8'b00100000 ;
56 :dout = 8'b00100010 ;
57 :dout = 8'b00011100 ;
67 :dout = 8'b00111100 ;
68 :dout = 8'b00010010 ;
69 :dout = 8'b00010010 ;
70 :dout = 8'b00010010 ;
71 :dout = 8'b00010010 ;
72 :dout = 8'b00010010 ;
73 :dout = 8'b00111100 ;
83 :dout = 8'b00111110 ;
84 :dout = 8'b00100000 ;
85 :dout = 8'b00100000 ;
86 :dout = 8'b00111000 ;
87 :dout = 8'b00100000 ;
88 :dout = 8'b00100000 ;
89 :dout = 8'b00111110 ;
99 :dout = 8'b00111110 ;
100 :dout = 8'b00100000 ;
101 :dout = 8'b00100000 ;
102 :dout = 8'b00111100 ;
103 :dout = 8'b00100000 ;
104 :dout = 8'b00100000 ;
105 :dout = 8'b00100000 ;
115 :dout = 8'b00011110 ;
116 :dout = 8'b00100000 ;
117 :dout = 8'b00100000 ;
118 :dout = 8'b00100110 ;
119 :dout = 8'b00100010 ;
120 :dout = 8'b00100010 ;
121 :dout = 8'b00011110 ;
131 :dout = 8'b00100010 ;
132 :dout = 8'b00100010 ;
133 :dout = 8'b00100010 ;
134 :dout = 8'b00111110 ;
135 :dout = 8'b00100010 ;
136 :dout = 8'b00100010 ;
137 :dout = 8'b00100010 ;
147 :dout = 8'b00011100 ;
148 :dout = 8'b00001000 ;
149 :dout = 8'b00001000 ;
150 :dout = 8'b00001000 ;
151 :dout = 8'b00001000 ;
152 :dout = 8'b00001000 ;
153 :dout = 8'b00011100 ;
163 :dout = 8'b00000010 ;
164 :dout = 8'b00000010 ;
165 :dout = 8'b00000010 ;
166 :dout = 8'b00000010 ;
167 :dout = 8'b00100010 ;
168 :dout = 8'b00100010 ;
169 :dout = 8'b00011100 ;
179 :dout = 8'b00100010 ;
180 :dout = 8'b00100100 ;
181 :dout = 8'b00101000 ;
182 :dout = 8'b00110000 ;
183 :dout = 8'b00110000 ;
184 :dout = 8'b00101000 ;
185 :dout = 8'b00100100 ;
195 :dout = 8'b00100000 ;
196 :dout = 8'b00100000 ;
197 :dout = 8'b00100000 ;
198 :dout = 8'b00100000 ;
199 :dout = 8'b00100000 ;
200 :dout = 8'b00100000 ;
201 :dout = 8'b00111110 ;
211 :dout = 8'b00100010 ;
212 :dout = 8'b00110110 ;
213 :dout = 8'b00101010 ;
214 :dout = 8'b00100010 ;
215 :dout = 8'b00100010 ;
216 :dout = 8'b00100010 ;
217 :dout = 8'b00100010 ;
227 :dout = 8'b00100010 ;
228 :dout = 8'b00110010 ;
229 :dout = 8'b00101010 ;
230 :dout = 8'b00100110 ;
231 :dout = 8'b00100010 ;
232 :dout = 8'b00100010 ;
233 :dout = 8'b00100010 ;
243 :dout = 8'b00011100 ;
244 :dout = 8'b00100010 ;
245 :dout = 8'b00100010 ;
246 :dout = 8'b00100010 ;
247 :dout = 8'b00100010 ;
248 :dout = 8'b00100010 ;
249 :dout = 8'b00011100 ;
259 :dout = 8'b00111100 ;
260 :dout = 8'b00100010 ;
261 :dout = 8'b00100010 ;
262 :dout = 8'b00111100 ;
263 :dout = 8'b00100000 ;
264 :dout = 8'b00100000 ;
265 :dout = 8'b00100000 ;
275 :dout = 8'b00011100 ;
276 :dout = 8'b00100010 ;
277 :dout = 8'b00100010 ;
278 :dout = 8'b00100010 ;
279 :dout = 8'b00101010 ;
280 :dout = 8'b00100100 ;
281 :dout = 8'b00011010 ;
291 :dout = 8'b00111100 ;
292 :dout = 8'b00100010 ;
293 :dout = 8'b00100010 ;
294 :dout = 8'b00111100 ;
295 :dout = 8'b00101000 ;
296 :dout = 8'b00100100 ;
297 :dout = 8'b00100010 ;
307 :dout = 8'b00011100 ;
308 :dout = 8'b00100010 ;
309 :dout = 8'b00010000 ;
310 :dout = 8'b00001000 ;
311 :dout = 8'b00000100 ;
312 :dout = 8'b00100010 ;
313 :dout = 8'b00011100 ;
323 :dout = 8'b00111110 ;
324 :dout = 8'b00001000 ;
325 :dout = 8'b00001000 ;
326 :dout = 8'b00001000 ;
327 :dout = 8'b00001000 ;
328 :dout = 8'b00001000 ;
329 :dout = 8'b00001000 ;
339 :dout = 8'b00100010 ;
340 :dout = 8'b00100010 ;
341 :dout = 8'b00100010 ;
342 :dout = 8'b00100010 ;
343 :dout = 8'b00100010 ;
344 :dout = 8'b00100010 ;
345 :dout = 8'b00011100 ;
355 :dout = 8'b00100010 ;
356 :dout = 8'b00100010 ;
357 :dout = 8'b00100010 ;
358 :dout = 8'b00100010 ;
359 :dout = 8'b00010100 ;
360 :dout = 8'b00010100 ;
361 :dout = 8'b00001000 ;
371 :dout = 8'b00100010 ;
372 :dout = 8'b00100010 ;
373 :dout = 8'b00100010 ;
374 :dout = 8'b00100010 ;
375 :dout = 8'b00101010 ;
376 :dout = 8'b00110110 ;
377 :dout = 8'b00100010 ;
387 :dout = 8'b00100010 ;
388 :dout = 8'b00100010 ;
389 :dout = 8'b00010100 ;
390 :dout = 8'b00001000 ;
391 :dout = 8'b00010100 ;
392 :dout = 8'b00100010 ;
393 :dout = 8'b00100010 ;
403 :dout = 8'b00100010 ;
404 :dout = 8'b00100010 ;
405 :dout = 8'b00010100 ;
406 :dout = 8'b00001000 ;
407 :dout = 8'b00001000 ;
408 :dout = 8'b00001000 ;
409 :dout = 8'b00001000 ;
419 :dout = 8'b00111110 ;
420 :dout = 8'b00000010 ;
421 :dout = 8'b00000100 ;
422 :dout = 8'b00001000 ;
423 :dout = 8'b00010000 ;
424 :dout = 8'b00100000 ;
425 :dout = 8'b00111110 ;
435 :dout = 8'b00011100 ;
436 :dout = 8'b00010000 ;
437 :dout = 8'b00010000 ;
438 :dout = 8'b00010000 ;
439 :dout = 8'b00010000 ;
440 :dout = 8'b00010000 ;
441 :dout = 8'b00011100 ;
451 :dout = 8'b00100000 ;
452 :dout = 8'b00100000 ;
453 :dout = 8'b00010000 ;
454 :dout = 8'b00001000 ;
455 :dout = 8'b00000100 ;
456 :dout = 8'b00000010 ;
457 :dout = 8'b00000010 ;
467 :dout = 8'b00011100 ;
468 :dout = 8'b00000100 ;
469 :dout = 8'b00000100 ;
470 :dout = 8'b00000100 ;
471 :dout = 8'b00000100 ;
472 :dout = 8'b00000100 ;
473 :dout = 8'b00011100 ;
483 :dout = 8'b00001000 ;
484 :dout = 8'b00011100 ;
485 :dout = 8'b00111110 ;
486 :dout = 8'b00001000 ;
487 :dout = 8'b00001000 ;
488 :dout = 8'b00001000 ;
489 :dout = 8'b00001000 ;
500 :dout = 8'b00001000 ;
501 :dout = 8'b00010000 ;
502 :dout = 8'b00111110 ;
503 :dout = 8'b00010000 ;
504 :dout = 8'b00001000 ;
531 :dout = 8'b00001000 ;
532 :dout = 8'b00001000 ;
533 :dout = 8'b00001000 ;
534 :dout = 8'b00001000 ;
535 :dout = 8'b00001000 ;
537 :dout = 8'b00001000 ;
547 :dout = 8'b00010100 ;
548 :dout = 8'b00010100 ;
563 :dout = 8'b00010100 ;
564 :dout = 8'b00010100 ;
565 :dout = 8'b00110110 ;
567 :dout = 8'b00110110 ;
568 :dout = 8'b00010100 ;
569 :dout = 8'b00010100 ;
579 :dout = 8'b00001000 ;
580 :dout = 8'b00011110 ;
581 :dout = 8'b00100000 ;
582 :dout = 8'b00011100 ;
583 :dout = 8'b00000010 ;
584 :dout = 8'b00111100 ;
585 :dout = 8'b00001000 ;
595 :dout = 8'b00110010 ;
596 :dout = 8'b00110010 ;
597 :dout = 8'b00000100 ;
598 :dout = 8'b00001000 ;
599 :dout = 8'b00010000 ;
600 :dout = 8'b00100110 ;
601 :dout = 8'b00100110 ;
611 :dout = 8'b00010000 ;
612 :dout = 8'b00101000 ;
613 :dout = 8'b00101000 ;
614 :dout = 8'b00010010 ;
615 :dout = 8'b00101100 ;
616 :dout = 8'b00101100 ;
617 :dout = 8'b00010010 ;
627 :dout = 8'b00001000 ;
628 :dout = 8'b00001000 ;
643 :dout = 8'b00000100 ;
644 :dout = 8'b00001000 ;
645 :dout = 8'b00010000 ;
646 :dout = 8'b00010000 ;
647 :dout = 8'b00010000 ;
648 :dout = 8'b00001000 ;
649 :dout = 8'b00000100 ;
659 :dout = 8'b00010000 ;
660 :dout = 8'b00001000 ;
661 :dout = 8'b00000100 ;
662 :dout = 8'b00000100 ;
663 :dout = 8'b00000100 ;
664 :dout = 8'b00001000 ;
665 :dout = 8'b00010000 ;
676 :dout = 8'b00001000 ;
677 :dout = 8'b00101010 ;
678 :dout = 8'b00011100 ;
679 :dout = 8'b00101010 ;
680 :dout = 8'b00001000 ;
692 :dout = 8'b00001000 ;
693 :dout = 8'b00001000 ;
694 :dout = 8'b00111110 ;
695 :dout = 8'b00001000 ;
696 :dout = 8'b00001000 ;
710 :dout = 8'b00001100 ;
711 :dout = 8'b00001100 ;
712 :dout = 8'b00000100 ;
713 :dout = 8'b00001000 ;
726 :dout = 8'b00111110 ;
744 :dout = 8'b00001000 ;
745 :dout = 8'b00001000 ;
755 :dout = 8'b00000010 ;
756 :dout = 8'b00000010 ;
757 :dout = 8'b00000100 ;
758 :dout = 8'b00001000 ;
759 :dout = 8'b00010000 ;
760 :dout = 8'b00100000 ;
761 :dout = 8'b00100000 ;
771 :dout = 8'b00011100 ;
772 :dout = 8'b00100010 ;
773 :dout = 8'b00100110 ;
774 :dout = 8'b00101010 ;
775 :dout = 8'b00110010 ;
776 :dout = 8'b00100010 ;
777 :dout = 8'b00011100 ;
787 :dout = 8'b00001000 ;
788 :dout = 8'b00011000 ;
789 :dout = 8'b00001000 ;
790 :dout = 8'b00001000 ;
791 :dout = 8'b00001000 ;
792 :dout = 8'b00001000 ;
793 :dout = 8'b00011100 ;
803 :dout = 8'b00011100 ;
804 :dout = 8'b00100010 ;
805 :dout = 8'b00000010 ;
806 :dout = 8'b00011100 ;
807 :dout = 8'b00100000 ;
808 :dout = 8'b00100000 ;
809 :dout = 8'b00111110 ;
819 :dout = 8'b00011100 ;
820 :dout = 8'b00100010 ;
821 :dout = 8'b00000010 ;
822 :dout = 8'b00001100 ;
823 :dout = 8'b00000010 ;
824 :dout = 8'b00100010 ;
825 :dout = 8'b00011100 ;
835 :dout = 8'b00000100 ;
836 :dout = 8'b00001100 ;
837 :dout = 8'b00010100 ;
838 :dout = 8'b00111110 ;
839 :dout = 8'b00000100 ;
840 :dout = 8'b00000100 ;
841 :dout = 8'b00000100 ;
851 :dout = 8'b00111110 ;
852 :dout = 8'b00100000 ;
853 :dout = 8'b00111100 ;
854 :dout = 8'b00000010 ;
855 :dout = 8'b00000010 ;
856 :dout = 8'b00100010 ;
857 :dout = 8'b00011100 ;
867 :dout = 8'b00011100 ;
868 :dout = 8'b00100000 ;
869 :dout = 8'b00100000 ;
870 :dout = 8'b00111100 ;
871 :dout = 8'b00100010 ;
872 :dout = 8'b00100010 ;
873 :dout = 8'b00011100 ;
883 :dout = 8'b00111110 ;
884 :dout = 8'b00000010 ;
885 :dout = 8'b00000100 ;
886 :dout = 8'b00001000 ;
887 :dout = 8'b00010000 ;
888 :dout = 8'b00100000 ;
889 :dout = 8'b00100000 ;
899 :dout = 8'b00011100 ;
900 :dout = 8'b00100010 ;
901 :dout = 8'b00100010 ;
902 :dout = 8'b00011100 ;
903 :dout = 8'b00100010 ;
904 :dout = 8'b00100010 ;
905 :dout = 8'b00011100 ;
915 :dout = 8'b00011100 ;
916 :dout = 8'b00100010 ;
917 :dout = 8'b00100010 ;
918 :dout = 8'b00011110 ;
919 :dout = 8'b00000010 ;
920 :dout = 8'b00000010 ;
921 :dout = 8'b00011100 ;
933 :dout = 8'b00001000 ;
935 :dout = 8'b00001000 ;
947 :dout = 8'b00001100 ;
948 :dout = 8'b00001100 ;
950 :dout = 8'b00001100 ;
951 :dout = 8'b00001100 ;
952 :dout = 8'b00000100 ;
953 :dout = 8'b00001000 ;
963 :dout = 8'b00000100 ;
964 :dout = 8'b00001000 ;
965 :dout = 8'b00010000 ;
966 :dout = 8'b00100000 ;
967 :dout = 8'b00010000 ;
968 :dout = 8'b00001000 ;
969 :dout = 8'b00000100 ;
981 :dout = 8'b00111110 ;
983 :dout = 8'b00111110 ;
995 :dout = 8'b00100000 ;
996 :dout = 8'b00010000 ;
997 :dout = 8'b00001000 ;
998 :dout = 8'b00000100 ;
999 :dout = 8'b00001000 ;
1000 :dout = 8'b00010000 ;
1001 :dout = 8'b00100000 ;
1011 :dout = 8'b00011100 ;
1012 :dout = 8'b00100010 ;
1013 :dout = 8'b00000100 ;
1014 :dout = 8'b00001000 ;
1015 :dout = 8'b00001000 ;
1017 :dout = 8'b00001000 ;
default :dout = 8'b00000000 ;
endcase
end

endmodule


